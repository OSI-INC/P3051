---------- RING OSCILLATOR ENTITY DECLARATION ----------
library ieee;  
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ring_oscillator is 
	generic (
		ring_len : integer := 15);
	port (
		ENABLE : in std_logic;
		CK : out std_logic);
end;

architecture behavior of ring_oscillator is 

-- Unlike previous versions of our ring oscillator, this one operates on a 
-- a simple principle: keep adding gates to the ring until you get the correct
-- period. The trick is to avoid consuming power with gates that we don't 
-- use. So long as we use all the gates in the ring, the current consumpiont
-- of the ring is independent of the number of gates, but as soon as we start
-- running unused gates off the ring, these will consume power.

-- When compiling and routing this oscillator, we have to convince the VHDL 
-- compiler to retain the ring buffers, despite its great desire to elimnate 
-- them all, and its complaints that we have timing loops. In a LCMXO2-1200ZE 
-- with core power supply dropped to 1.0 V, the gate delay is around 3.5 ns. 
-- For each gate we add to the ring oscillator, we increase the period by 
-- roughly 7.0 ns, which is ample resolution for the generation of a period 
-- in the range 195-215 ns. 

-- Functions and Procedures	
	function to_std_logic (v: boolean) return std_ulogic is
	begin if v then return('1'); else return('0'); end if; end function;

-- Attributes to guide the compiler.
	attribute syn_keep : boolean;
	attribute nomerge : string;

-- Ring Oscillator and Transmit Clock
	component BUFBA is port (A : in std_logic; Z : out std_logic); end component;
	signal R : std_logic_vector(ring_len downto 0);
	attribute syn_keep of R : signal is true;
	attribute nomerge of R : signal is ""; 

begin

-- Declare the ring oscillator gate entities.
	gen_ring : for i in 0 to ring_len-1 generate
        stage : BUFBA
            port map (
                A => R(i),
                Z => R(i+1)
            );
    end generate;

-- When ENABLE, feed back the output of the final gate to the first gate.
	R(0) <= to_std_logic((ENABLE = '1') and (R(ring_len) = '0'));
	
-- The clock output.
	CK <= R(0);
end behavior;
------------ END RING OSCILLATOR DECLARATION -----------


----------- POWER CONTROL UNIT ENTITY DECLARATION ------
-- VHDL netlist generated by SCUBA Diamond_2.2_Production (99)
-- Tue Aug 19 11:48:15 2014

library IEEE;
use IEEE.std_logic_1164.all;
-- synopsys translate_off
library MACHXO2;
use MACHXO2.components.all;
-- synopsys translate_on

entity PCU is
    port (
        USERSTDBY: in  std_logic; 
        CLRFLAG: in  std_logic; 
        STDBY: out  std_logic; 
        SFLAG: out  std_logic);
end PCU;

architecture Structure of PCU is

    -- internal signal declarations
    signal scuba_vlo: std_logic;

    -- local component declarations
    component VLO
        port (Z: out  std_logic);
    end component;
    component PCNTR
        generic (STDBYOPT : in String; TIMEOUT : in String; 
                WAKEUP : in String; POROFF : in String; 
                BGOFF : in String);
        port (CLK: in  std_logic; USERTIMEOUT: in  std_logic; 
            USERSTDBY: in  std_logic; CLRFLAG: in  std_logic; 
            CFGWAKE: in  std_logic; CFGSTDBY: in  std_logic; 
            STDBY: out  std_logic; STOP: out  std_logic; 
            SFLAG: out  std_logic);
    end component;
    attribute NGD_DRC_MASK : integer;
    attribute NGD_DRC_MASK of Structure : architecture is 1;

begin
    -- component instantiation statements
    scuba_vlo_inst: VLO
        port map (Z=>scuba_vlo);

    PCNTR_Inst0: PCNTR
        generic map (BGOFF=> "TRUE", POROFF=> "TRUE", WAKEUP=> "USER", 
        TIMEOUT=> "BYPASS", STDBYOPT=> "USER")
        port map (CLK=>scuba_vlo, USERTIMEOUT=>scuba_vlo, 
            USERSTDBY=>USERSTDBY, CLRFLAG=>CLRFLAG, CFGWAKE=>scuba_vlo, 
            CFGSTDBY=>scuba_vlo, STDBY=>STDBY, STOP=>open, SFLAG=>SFLAG);

end Structure;
----------- END POWER CONTROL UNIT ENTITY DECLARATION ------
