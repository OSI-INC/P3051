---------- RING OSCILLATOR ENTITY DECLARATION ----------
library ieee;  
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ring_oscillator is 
	generic (
		calib_range : integer := 15);
	port (
		ENABLE : in std_logic;
		calib : in integer range 0 to calib_range;
		CK : out std_logic);
end;

architecture behavior of ring_oscillator is 

-- WARNING: The ring oscillator is precarious, in that it is hard to predict what
-- small changes in the code will do to its behavior.

-- When compiling and routing this oscillator, we have to convince the VHDL compiler
-- to retain four buffers to make the ring, despite its great desire to elimnate them
-- all, and its complaints that we have timing loops. On the LCMXO2-1200ZE-1U, our 
-- four-gate ring runs at about 140 MHz, implying an individual gate delay of 0.8 ns. 
-- The compiler calculates there is no way the chip can count a 140-MHz clock in a 
-- 5-bit counter, so we don't tell it the true speed of the ring when we perform timing 
-- analysis. If we were to increase the ring to five gates, we would no longer have the 
-- resolution in CK period adjustment to guarantee that the period is within the 
-- 195-215 ns interval acceptable for SCT messages.

-- Functions and Procedures	
	function to_std_logic (v: boolean) return std_ulogic is
	begin if v then return('1'); else return('0'); end if; end function;

-- Attributes to guide the compiler.
	attribute syn_keep : boolean;
	attribute nomerge : string;

-- Ring Oscillator and Transmit Clock
	component BUFBA is port (A : in std_logic; Z : out std_logic); end component;
	signal RIN, R1, R2, R3, R4, R5, R6 : std_logic;
	attribute syn_keep of RIN, R1, R2, R3, R4, R5, R6 : signal is true;
	attribute nomerge of RIN, R1, R2, R3, R4, R5, R6 : signal is ""; 

begin

-- Declare the ring oscillator gate entities.
	ring1 : BUFBA port map (RIN,R1);
	ring2 : BUFBA port map (R1,R2);
	ring3 : BUFBA port map (R2,R3);
	ring4 : BUFBA port map (R3,R4);
	ring5 : BUFBA port map (R4,R5);
	ring6 : BUFBA port map (R5,R6);

-- When ENABLE, feed back the output of one of the gates to the first gate 
-- in the ring. The ring needs to oscillate fast enough that integer fractions
-- of the frequency will get us close to our ideal output frequency. It must
-- run slow enough that our dividor can function.
	RIN <= to_std_logic((ENABLE = '1') and (R3 = '0'));
	
-- The divider process takes the ring osillator output and divides it down to
-- a slower frequency. When the divisor is even, the output clock will have 
-- exactly 50% duty cycle. When odd, the duty cycle will be as close to 50% as
-- we can get.
	divider : process (RIN) is
		variable count, next_count : integer range 0 to calib_range;
	begin	
		
		-- Act on the rising edge of RIN.
		if rising_edge(RIN) then
		
			-- Count down from calib to zero, a total of calib+1 RIN periods
			-- will make up the output clock period.
			if (count = 0) then 
				next_count := calib;
			else 
				next_count := count - 1;
			end if;
			
			-- We try to get close to 50% duty cycle. We don't use feedback,
			-- but instead specify fully the values of CK in terms of calib 
			-- for all values of count so as to speed up the logic behind CK. 
			if (count <= calib/2) then
				CK <= '1';
			else
				CK <= '0';
			end if;
			
			-- Se the next count.
			count := next_count;
		end if;
	end process;
end behavior;
------------ END RING OSCILLATOR DECLARATION -----------


----------- POWER CONTROL UNIT ENTITY DECLARATION ------
-- VHDL netlist generated by SCUBA Diamond_2.2_Production (99)
-- Tue Aug 19 11:48:15 2014

library IEEE;
use IEEE.std_logic_1164.all;
-- synopsys translate_off
library MACHXO2;
use MACHXO2.components.all;
-- synopsys translate_on

entity PCU is
    port (
        USERSTDBY: in  std_logic; 
        CLRFLAG: in  std_logic; 
        STDBY: out  std_logic; 
        SFLAG: out  std_logic);
end PCU;

architecture Structure of PCU is

    -- internal signal declarations
    signal scuba_vlo: std_logic;

    -- local component declarations
    component VLO
        port (Z: out  std_logic);
    end component;
    component PCNTR
        generic (STDBYOPT : in String; TIMEOUT : in String; 
                WAKEUP : in String; POROFF : in String; 
                BGOFF : in String);
        port (CLK: in  std_logic; USERTIMEOUT: in  std_logic; 
            USERSTDBY: in  std_logic; CLRFLAG: in  std_logic; 
            CFGWAKE: in  std_logic; CFGSTDBY: in  std_logic; 
            STDBY: out  std_logic; STOP: out  std_logic; 
            SFLAG: out  std_logic);
    end component;
    attribute NGD_DRC_MASK : integer;
    attribute NGD_DRC_MASK of Structure : architecture is 1;

begin
    -- component instantiation statements
    scuba_vlo_inst: VLO
        port map (Z=>scuba_vlo);

    PCNTR_Inst0: PCNTR
        generic map (BGOFF=> "TRUE", POROFF=> "TRUE", WAKEUP=> "USER", 
        TIMEOUT=> "BYPASS", STDBYOPT=> "USER")
        port map (CLK=>scuba_vlo, USERTIMEOUT=>scuba_vlo, 
            USERSTDBY=>USERSTDBY, CLRFLAG=>CLRFLAG, CFGWAKE=>scuba_vlo, 
            CFGSTDBY=>scuba_vlo, STDBY=>STDBY, STOP=>open, SFLAG=>SFLAG);

end Structure;
----------- END POWER CONTROL UNIT ENTITY DECLARATION ------
